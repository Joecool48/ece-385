// final_project.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module final_project (
		input  wire        avalon_control_fixed_location,  //     avalon_control.fixed_location
		input  wire [31:0] avalon_control_read_base,       //                   .read_base
		input  wire [31:0] avalon_control_read_length,     //                   .read_length
		input  wire        avalon_control_go,              //                   .go
		output wire        avalon_control_done,            //                   .done
		output wire        avalon_control_early_done,      //                   .early_done
		input  wire        avalon_user_read_buffer,        //        avalon_user.read_buffer
		output wire [7:0]  avalon_user_buffer_output_data, //                   .buffer_output_data
		output wire        avalon_user_data_available,     //                   .data_available
		input  wire        clk_clk,                        //                clk.clk
		input  wire        reset_reset_n,                  //              reset.reset_n
		output wire        sdram_clk_clk,                  //          sdram_clk.clk
		output wire [11:0] sdram_wire_addr,                //         sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                  //                   .ba
		output wire        sdram_wire_cas_n,               //                   .cas_n
		output wire        sdram_wire_cke,                 //                   .cke
		output wire        sdram_wire_cs_n,                //                   .cs_n
		inout  wire [31:0] sdram_wire_dq,                  //                   .dq
		output wire [3:0]  sdram_wire_dqm,                 //                   .dqm
		output wire        sdram_wire_ras_n,               //                   .ras_n
		output wire        sdram_wire_we_n,                //                   .we_n
		output wire [31:0] sprite_address_pio_export,      // sprite_address_pio.export
		output wire [15:0] sprite_height_pio_export,       //  sprite_height_pio.export
		output wire [15:0] sprite_id_pio_export,           //      sprite_id_pio.export
		output wire [15:0] sprite_width_pio_export,        //   sprite_width_pio.export
		output wire [15:0] sprite_x_pio_export,            //       sprite_x_pio.export
		output wire [15:0] sprite_y_pio_export,            //       sprite_y_pio.export
		output wire        sys_clk_clk                     //            sys_clk.clk
	);

	wire         pll_c0_clk;                                                     // pll:c0 -> [irq_mapper:clk, jtag_game_nios:clk, master_template_0:clk, mm_interconnect_0:pll_c0_clk, nios2_gen2_0:clk, rst_controller:clk, sdram:clk, sprite_address_pio:clk, sprite_height_pio:clk, sprite_id_pio:clk, sprite_width_pio:clk, sprite_x_pio:clk, sprite_y_pio:clk, sysid:clock]
	wire   [7:0] master_template_0_avalon_master_readdata;                       // mm_interconnect_0:master_template_0_avalon_master_readdata -> master_template_0:master_readdata
	wire         master_template_0_avalon_master_waitrequest;                    // mm_interconnect_0:master_template_0_avalon_master_waitrequest -> master_template_0:master_waitrequest
	wire  [31:0] master_template_0_avalon_master_address;                        // master_template_0:master_address -> mm_interconnect_0:master_template_0_avalon_master_address
	wire         master_template_0_avalon_master_read;                           // master_template_0:master_read -> mm_interconnect_0:master_template_0_avalon_master_read
	wire         master_template_0_avalon_master_byteenable;                     // master_template_0:master_byteenable -> mm_interconnect_0:master_template_0_avalon_master_byteenable
	wire         master_template_0_avalon_master_readdatavalid;                  // mm_interconnect_0:master_template_0_avalon_master_readdatavalid -> master_template_0:master_readdatavalid
	wire   [6:0] master_template_0_avalon_master_burstcount;                     // master_template_0:master_burstcount -> mm_interconnect_0:master_template_0_avalon_master_burstcount
	wire  [31:0] nios2_gen2_0_data_master_readdata;                              // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                           // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                           // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [24:0] nios2_gen2_0_data_master_address;                               // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                            // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                  // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                                 // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                             // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                       // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [24:0] nios2_gen2_0_instruction_master_address;                        // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                           // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_chipselect -> jtag_game_nios:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_readdata;    // jtag_game_nios:av_readdata -> mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_waitrequest; // jtag_game_nios:av_waitrequest -> mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_address -> jtag_game_nios:av_address
	wire         mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_read -> jtag_game_nios:av_read_n
	wire         mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_write -> jtag_game_nios:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_game_nios_avalon_jtag_slave_writedata -> jtag_game_nios:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                 // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                  // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;        // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;     // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;     // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;       // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                          // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                            // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                         // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                             // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                          // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                       // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                               // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                           // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                       // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                        // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                           // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                          // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                      // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_sprite_id_pio_s1_chipselect;                  // mm_interconnect_0:sprite_id_pio_s1_chipselect -> sprite_id_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_id_pio_s1_readdata;                    // sprite_id_pio:readdata -> mm_interconnect_0:sprite_id_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_id_pio_s1_address;                     // mm_interconnect_0:sprite_id_pio_s1_address -> sprite_id_pio:address
	wire         mm_interconnect_0_sprite_id_pio_s1_write;                       // mm_interconnect_0:sprite_id_pio_s1_write -> sprite_id_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_id_pio_s1_writedata;                   // mm_interconnect_0:sprite_id_pio_s1_writedata -> sprite_id_pio:writedata
	wire         mm_interconnect_0_sprite_address_pio_s1_chipselect;             // mm_interconnect_0:sprite_address_pio_s1_chipselect -> sprite_address_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_address_pio_s1_readdata;               // sprite_address_pio:readdata -> mm_interconnect_0:sprite_address_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_address_pio_s1_address;                // mm_interconnect_0:sprite_address_pio_s1_address -> sprite_address_pio:address
	wire         mm_interconnect_0_sprite_address_pio_s1_write;                  // mm_interconnect_0:sprite_address_pio_s1_write -> sprite_address_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_address_pio_s1_writedata;              // mm_interconnect_0:sprite_address_pio_s1_writedata -> sprite_address_pio:writedata
	wire         mm_interconnect_0_sprite_width_pio_s1_chipselect;               // mm_interconnect_0:sprite_width_pio_s1_chipselect -> sprite_width_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_width_pio_s1_readdata;                 // sprite_width_pio:readdata -> mm_interconnect_0:sprite_width_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_width_pio_s1_address;                  // mm_interconnect_0:sprite_width_pio_s1_address -> sprite_width_pio:address
	wire         mm_interconnect_0_sprite_width_pio_s1_write;                    // mm_interconnect_0:sprite_width_pio_s1_write -> sprite_width_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_width_pio_s1_writedata;                // mm_interconnect_0:sprite_width_pio_s1_writedata -> sprite_width_pio:writedata
	wire         mm_interconnect_0_sprite_height_pio_s1_chipselect;              // mm_interconnect_0:sprite_height_pio_s1_chipselect -> sprite_height_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_height_pio_s1_readdata;                // sprite_height_pio:readdata -> mm_interconnect_0:sprite_height_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_height_pio_s1_address;                 // mm_interconnect_0:sprite_height_pio_s1_address -> sprite_height_pio:address
	wire         mm_interconnect_0_sprite_height_pio_s1_write;                   // mm_interconnect_0:sprite_height_pio_s1_write -> sprite_height_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_height_pio_s1_writedata;               // mm_interconnect_0:sprite_height_pio_s1_writedata -> sprite_height_pio:writedata
	wire         mm_interconnect_0_sprite_x_pio_s1_chipselect;                   // mm_interconnect_0:sprite_x_pio_s1_chipselect -> sprite_x_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_x_pio_s1_readdata;                     // sprite_x_pio:readdata -> mm_interconnect_0:sprite_x_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_x_pio_s1_address;                      // mm_interconnect_0:sprite_x_pio_s1_address -> sprite_x_pio:address
	wire         mm_interconnect_0_sprite_x_pio_s1_write;                        // mm_interconnect_0:sprite_x_pio_s1_write -> sprite_x_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_x_pio_s1_writedata;                    // mm_interconnect_0:sprite_x_pio_s1_writedata -> sprite_x_pio:writedata
	wire         mm_interconnect_0_sprite_y_pio_s1_chipselect;                   // mm_interconnect_0:sprite_y_pio_s1_chipselect -> sprite_y_pio:chipselect
	wire  [31:0] mm_interconnect_0_sprite_y_pio_s1_readdata;                     // sprite_y_pio:readdata -> mm_interconnect_0:sprite_y_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_sprite_y_pio_s1_address;                      // mm_interconnect_0:sprite_y_pio_s1_address -> sprite_y_pio:address
	wire         mm_interconnect_0_sprite_y_pio_s1_write;                        // mm_interconnect_0:sprite_y_pio_s1_write -> sprite_y_pio:write_n
	wire  [31:0] mm_interconnect_0_sprite_y_pio_s1_writedata;                    // mm_interconnect_0:sprite_y_pio_s1_writedata -> sprite_y_pio:writedata
	wire         irq_mapper_receiver0_irq;                                       // jtag_game_nios:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                           // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [irq_mapper:reset, jtag_game_nios:rst_n, master_template_0:reset, mm_interconnect_0:master_template_0_clock_reset_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, sdram:reset_n, sprite_address_pio:reset_n, sprite_height_pio:reset_n, sprite_id_pio:reset_n, sprite_width_pio:reset_n, sprite_x_pio:reset_n, sprite_y_pio:reset_n, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	final_project_jtag_game_nios jtag_game_nios (
		.clk            (pll_c0_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                        //               irq.irq
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (8),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (1),
		.MAXIMUM_BURST_COUNT (64),
		.BURST_COUNT_WIDTH   (7),
		.FIFO_DEPTH          (128),
		.FIFO_DEPTH_LOG2     (7),
		.MEMORY_BASED_FIFO   (1)
	) master_template_0 (
		.clk                     (pll_c0_clk),                                    //       clock_reset.clk
		.reset                   (rst_controller_reset_out_reset),                // clock_reset_reset.reset
		.master_address          (master_template_0_avalon_master_address),       //     avalon_master.address
		.master_read             (master_template_0_avalon_master_read),          //                  .read
		.master_byteenable       (master_template_0_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (master_template_0_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (master_template_0_avalon_master_readdatavalid), //                  .readdatavalid
		.master_burstcount       (master_template_0_avalon_master_burstcount),    //                  .burstcount
		.master_waitrequest      (master_template_0_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (avalon_control_fixed_location),                 //           control.export
		.control_read_base       (avalon_control_read_base),                      //                  .export
		.control_read_length     (avalon_control_read_length),                    //                  .export
		.control_go              (avalon_control_go),                             //                  .export
		.control_done            (avalon_control_done),                           //                  .export
		.control_early_done      (avalon_control_early_done),                     //                  .export
		.user_read_buffer        (avalon_user_read_buffer),                       //              user.export
		.user_buffer_output_data (avalon_user_buffer_output_data),                //                  .export
		.user_data_available     (avalon_user_data_available),                    //                  .export
		.master_write            (),                                              //       (terminated)
		.master_writedata        (),                                              //       (terminated)
		.control_write_base      (32'b00000000000000000000000000000000),          //       (terminated)
		.control_write_length    (32'b00000000000000000000000000000000),          //       (terminated)
		.user_write_buffer       (1'b0),                                          //       (terminated)
		.user_buffer_input_data  (8'b00000000),                                   //       (terminated)
		.user_buffer_full        ()                                               //       (terminated)
	);

	final_project_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (pll_c0_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                           //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	final_project_pll pll (
		.clk                (clk_clk),                                   //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0                 (pll_c0_clk),                                //                    c0.clk
		.c1                 (),                                          //                    c1.clk
		.c2                 (sdram_clk_clk),                             //                    c2.clk
		.c3                 (sys_clk_clk),                               //                    c3.clk
		.scandone           (),                                          //           (terminated)
		.scandataout        (),                                          //           (terminated)
		.areset             (1'b0),                                      //           (terminated)
		.locked             (),                                          //           (terminated)
		.phasedone          (),                                          //           (terminated)
		.phasecounterselect (4'b0000),                                   //           (terminated)
		.phaseupdown        (1'b0),                                      //           (terminated)
		.phasestep          (1'b0),                                      //           (terminated)
		.scanclk            (1'b0),                                      //           (terminated)
		.scanclkena         (1'b0),                                      //           (terminated)
		.scandata           (1'b0),                                      //           (terminated)
		.configupdate       (1'b0)                                       //           (terminated)
	);

	final_project_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_project_sprite_address_pio sprite_address_pio (
		.clk        (pll_c0_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (mm_interconnect_0_sprite_address_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_address_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_address_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_address_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_address_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_address_pio_export)                           // external_connection.export
	);

	final_project_sprite_height_pio sprite_height_pio (
		.clk        (pll_c0_clk),                                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_sprite_height_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_height_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_height_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_height_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_height_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_height_pio_export)                           // external_connection.export
	);

	final_project_sprite_height_pio sprite_id_pio (
		.clk        (pll_c0_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_sprite_id_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_id_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_id_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_id_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_id_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_id_pio_export)                           // external_connection.export
	);

	final_project_sprite_height_pio sprite_width_pio (
		.clk        (pll_c0_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_sprite_width_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_width_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_width_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_width_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_width_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_width_pio_export)                           // external_connection.export
	);

	final_project_sprite_height_pio sprite_x_pio (
		.clk        (pll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sprite_x_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_x_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_x_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_x_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_x_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_x_pio_export)                           // external_connection.export
	);

	final_project_sprite_height_pio sprite_y_pio (
		.clk        (pll_c0_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sprite_y_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sprite_y_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sprite_y_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sprite_y_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sprite_y_pio_s1_readdata),   //                    .readdata
		.out_port   (sprite_y_pio_export)                           // external_connection.export
	);

	final_project_sysid sysid (
		.clock    (pll_c0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	final_project_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                   (clk_clk),                                                        //                                                 clk_0_clk.clk
		.pll_c0_clk                                                      (pll_c0_clk),                                                     //                                                    pll_c0.clk
		.master_template_0_clock_reset_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // master_template_0_clock_reset_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset           (rst_controller_001_reset_out_reset),                             //           pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.master_template_0_avalon_master_address                         (master_template_0_avalon_master_address),                        //                           master_template_0_avalon_master.address
		.master_template_0_avalon_master_waitrequest                     (master_template_0_avalon_master_waitrequest),                    //                                                          .waitrequest
		.master_template_0_avalon_master_burstcount                      (master_template_0_avalon_master_burstcount),                     //                                                          .burstcount
		.master_template_0_avalon_master_byteenable                      (master_template_0_avalon_master_byteenable),                     //                                                          .byteenable
		.master_template_0_avalon_master_read                            (master_template_0_avalon_master_read),                           //                                                          .read
		.master_template_0_avalon_master_readdata                        (master_template_0_avalon_master_readdata),                       //                                                          .readdata
		.master_template_0_avalon_master_readdatavalid                   (master_template_0_avalon_master_readdatavalid),                  //                                                          .readdatavalid
		.nios2_gen2_0_data_master_address                                (nios2_gen2_0_data_master_address),                               //                                  nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                            (nios2_gen2_0_data_master_waitrequest),                           //                                                          .waitrequest
		.nios2_gen2_0_data_master_byteenable                             (nios2_gen2_0_data_master_byteenable),                            //                                                          .byteenable
		.nios2_gen2_0_data_master_read                                   (nios2_gen2_0_data_master_read),                                  //                                                          .read
		.nios2_gen2_0_data_master_readdata                               (nios2_gen2_0_data_master_readdata),                              //                                                          .readdata
		.nios2_gen2_0_data_master_write                                  (nios2_gen2_0_data_master_write),                                 //                                                          .write
		.nios2_gen2_0_data_master_writedata                              (nios2_gen2_0_data_master_writedata),                             //                                                          .writedata
		.nios2_gen2_0_data_master_debugaccess                            (nios2_gen2_0_data_master_debugaccess),                           //                                                          .debugaccess
		.nios2_gen2_0_instruction_master_address                         (nios2_gen2_0_instruction_master_address),                        //                           nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                     (nios2_gen2_0_instruction_master_waitrequest),                    //                                                          .waitrequest
		.nios2_gen2_0_instruction_master_read                            (nios2_gen2_0_instruction_master_read),                           //                                                          .read
		.nios2_gen2_0_instruction_master_readdata                        (nios2_gen2_0_instruction_master_readdata),                       //                                                          .readdata
		.jtag_game_nios_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_address),     //                          jtag_game_nios_avalon_jtag_slave.address
		.jtag_game_nios_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_write),       //                                                          .write
		.jtag_game_nios_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_read),        //                                                          .read
		.jtag_game_nios_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_readdata),    //                                                          .readdata
		.jtag_game_nios_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_writedata),   //                                                          .writedata
		.jtag_game_nios_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_waitrequest), //                                                          .waitrequest
		.jtag_game_nios_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_game_nios_avalon_jtag_slave_chipselect),  //                                                          .chipselect
		.nios2_gen2_0_debug_mem_slave_address                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),         //                              nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),           //                                                          .write
		.nios2_gen2_0_debug_mem_slave_read                               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),            //                                                          .read
		.nios2_gen2_0_debug_mem_slave_readdata                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),        //                                                          .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),       //                                                          .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),      //                                                          .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),     //                                                          .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),     //                                                          .debugaccess
		.pll_pll_slave_address                                           (mm_interconnect_0_pll_pll_slave_address),                        //                                             pll_pll_slave.address
		.pll_pll_slave_write                                             (mm_interconnect_0_pll_pll_slave_write),                          //                                                          .write
		.pll_pll_slave_read                                              (mm_interconnect_0_pll_pll_slave_read),                           //                                                          .read
		.pll_pll_slave_readdata                                          (mm_interconnect_0_pll_pll_slave_readdata),                       //                                                          .readdata
		.pll_pll_slave_writedata                                         (mm_interconnect_0_pll_pll_slave_writedata),                      //                                                          .writedata
		.sdram_s1_address                                                (mm_interconnect_0_sdram_s1_address),                             //                                                  sdram_s1.address
		.sdram_s1_write                                                  (mm_interconnect_0_sdram_s1_write),                               //                                                          .write
		.sdram_s1_read                                                   (mm_interconnect_0_sdram_s1_read),                                //                                                          .read
		.sdram_s1_readdata                                               (mm_interconnect_0_sdram_s1_readdata),                            //                                                          .readdata
		.sdram_s1_writedata                                              (mm_interconnect_0_sdram_s1_writedata),                           //                                                          .writedata
		.sdram_s1_byteenable                                             (mm_interconnect_0_sdram_s1_byteenable),                          //                                                          .byteenable
		.sdram_s1_readdatavalid                                          (mm_interconnect_0_sdram_s1_readdatavalid),                       //                                                          .readdatavalid
		.sdram_s1_waitrequest                                            (mm_interconnect_0_sdram_s1_waitrequest),                         //                                                          .waitrequest
		.sdram_s1_chipselect                                             (mm_interconnect_0_sdram_s1_chipselect),                          //                                                          .chipselect
		.sprite_address_pio_s1_address                                   (mm_interconnect_0_sprite_address_pio_s1_address),                //                                     sprite_address_pio_s1.address
		.sprite_address_pio_s1_write                                     (mm_interconnect_0_sprite_address_pio_s1_write),                  //                                                          .write
		.sprite_address_pio_s1_readdata                                  (mm_interconnect_0_sprite_address_pio_s1_readdata),               //                                                          .readdata
		.sprite_address_pio_s1_writedata                                 (mm_interconnect_0_sprite_address_pio_s1_writedata),              //                                                          .writedata
		.sprite_address_pio_s1_chipselect                                (mm_interconnect_0_sprite_address_pio_s1_chipselect),             //                                                          .chipselect
		.sprite_height_pio_s1_address                                    (mm_interconnect_0_sprite_height_pio_s1_address),                 //                                      sprite_height_pio_s1.address
		.sprite_height_pio_s1_write                                      (mm_interconnect_0_sprite_height_pio_s1_write),                   //                                                          .write
		.sprite_height_pio_s1_readdata                                   (mm_interconnect_0_sprite_height_pio_s1_readdata),                //                                                          .readdata
		.sprite_height_pio_s1_writedata                                  (mm_interconnect_0_sprite_height_pio_s1_writedata),               //                                                          .writedata
		.sprite_height_pio_s1_chipselect                                 (mm_interconnect_0_sprite_height_pio_s1_chipselect),              //                                                          .chipselect
		.sprite_id_pio_s1_address                                        (mm_interconnect_0_sprite_id_pio_s1_address),                     //                                          sprite_id_pio_s1.address
		.sprite_id_pio_s1_write                                          (mm_interconnect_0_sprite_id_pio_s1_write),                       //                                                          .write
		.sprite_id_pio_s1_readdata                                       (mm_interconnect_0_sprite_id_pio_s1_readdata),                    //                                                          .readdata
		.sprite_id_pio_s1_writedata                                      (mm_interconnect_0_sprite_id_pio_s1_writedata),                   //                                                          .writedata
		.sprite_id_pio_s1_chipselect                                     (mm_interconnect_0_sprite_id_pio_s1_chipselect),                  //                                                          .chipselect
		.sprite_width_pio_s1_address                                     (mm_interconnect_0_sprite_width_pio_s1_address),                  //                                       sprite_width_pio_s1.address
		.sprite_width_pio_s1_write                                       (mm_interconnect_0_sprite_width_pio_s1_write),                    //                                                          .write
		.sprite_width_pio_s1_readdata                                    (mm_interconnect_0_sprite_width_pio_s1_readdata),                 //                                                          .readdata
		.sprite_width_pio_s1_writedata                                   (mm_interconnect_0_sprite_width_pio_s1_writedata),                //                                                          .writedata
		.sprite_width_pio_s1_chipselect                                  (mm_interconnect_0_sprite_width_pio_s1_chipselect),               //                                                          .chipselect
		.sprite_x_pio_s1_address                                         (mm_interconnect_0_sprite_x_pio_s1_address),                      //                                           sprite_x_pio_s1.address
		.sprite_x_pio_s1_write                                           (mm_interconnect_0_sprite_x_pio_s1_write),                        //                                                          .write
		.sprite_x_pio_s1_readdata                                        (mm_interconnect_0_sprite_x_pio_s1_readdata),                     //                                                          .readdata
		.sprite_x_pio_s1_writedata                                       (mm_interconnect_0_sprite_x_pio_s1_writedata),                    //                                                          .writedata
		.sprite_x_pio_s1_chipselect                                      (mm_interconnect_0_sprite_x_pio_s1_chipselect),                   //                                                          .chipselect
		.sprite_y_pio_s1_address                                         (mm_interconnect_0_sprite_y_pio_s1_address),                      //                                           sprite_y_pio_s1.address
		.sprite_y_pio_s1_write                                           (mm_interconnect_0_sprite_y_pio_s1_write),                        //                                                          .write
		.sprite_y_pio_s1_readdata                                        (mm_interconnect_0_sprite_y_pio_s1_readdata),                     //                                                          .readdata
		.sprite_y_pio_s1_writedata                                       (mm_interconnect_0_sprite_y_pio_s1_writedata),                    //                                                          .writedata
		.sprite_y_pio_s1_chipselect                                      (mm_interconnect_0_sprite_y_pio_s1_chipselect),                   //                                                          .chipselect
		.sysid_control_slave_address                                     (mm_interconnect_0_sysid_control_slave_address),                  //                                       sysid_control_slave.address
		.sysid_control_slave_readdata                                    (mm_interconnect_0_sysid_control_slave_readdata)                  //                                                          .readdata
	);

	final_project_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
