module sys_manager ();